-------------------------------------------------------------------------------
-- Title      : Frame checker
-- Project    : MEEP
-------------------------------------------------------------------------------
-- File        : frame_check.vhd
-- Author      : Francelly K. Cano Ladino; francelly.canoladino@bsc.es
-- Company     : Barcelona Supercomputing Center (BSC)
-- Created     : 19/01/2021 - 19:12:35
-- Last update : Mon Feb 15 13:03:35 2021
-- Synthesizer : <Name> <version>
-- FPGA        : Alveo U280
-------------------------------------------------------------------------------
-- Description:  This module will implement a Frame checker to test a loopback using Aurora 64B/66B full-duplex connection.
-- With this module, we can check the frames generated by Frame_gen that arrive from Aurora Channel (RX).
-- We used the mas pseudo data algorithm to generate the same random data as Fram_Gen, using a comparator to check both values.
-- If an error is found, there is a counter that will increment each time.
-- Signals:
--   USER_CLK: The user_clk INPUT signal is a BUFG output deriving its input from tx_out_clk (Transceivers).   
--   RESET: This INPUT  signal reset the frame checker module.
--/User Interface: RX interface
--   AXIS_UI_RX_TDATA:This input signal is the random data that come from the AXI4-stream interface
--   (Aurora Channel)
--   AXIS_UI_RX_TVALID:This input signal indicates that this modules is driving a valid transfer.
--   DATA_ERROR_COUNT:This counter indicates if the comparison was unsuccessful incrementing each time occur an unmatch.
-- Comments : <Extra comments if they were needed>
-------------------------------------------------------------------------------
-- Copyright (c) 2019 DDR/TICH
-------------------------------------------------------------------------------
-- Revisions  : 1.0
-- Date/Time                Version               Engineer
-- dd/mm/yyyy - hh:mm        1.0             francelly.canoladino@bsc.es
-- Comments   : <Highlight the modifications>
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;
use ieee.STD_LOGIC_1164.all;
use ieee.std_logic_textio.all;
use std.textio.all;
use ieee.numeric_std.all;

entity frame_check is
  generic (

    DATA_WIDTH : integer := 64;
    STRB_WIDTH : integer := 8 -- STROBE bus width
    );
  port (

    -------------------------------------------------------------------------------
    -- System Interface
    -------------------------------------------------------------------------------     

    USER_CLK : in std_logic;            -- Aurora User Clk 
    RESET    : in std_logic;


    -------------------------------------------------------------------------------
    -- USER INTERFACE : RX INTERFACE
    -------------------------------------------------------------------------------

    AXIS_UI_RX_TDATA  : in  std_logic_vector(63 downto 0);
    AXIS_UI_RX_TVALID : in  std_logic;  --Handshake signal  
    DATA_ERR_COUNT    : out std_logic_vector(7 downto 0)

    );

end entity frame_check;

architecture rtl of frame_check is

-----------------------------------------------------------------------------
  -- CONSTANTS
-----------------------------------------------------------------------------
  constant AURORA_LANES     : integer                                      := 1;
  constant LANE_DATA_WIDTH  : integer                                      := (AURORA_LANES*64);
  constant REM_BUS          : integer                                      := 3;
-----------------------------------------------------------------------------
-- SIGNALS
-----------------------------------------------------------------------------
  signal reset_i            : std_logic                                    := '0';
  signal AXIS_UI_RX_TDATA_i : std_logic_vector(0 to (DATA_WIDTH-1))        := X"0000000000000000";
  signal r_rx_data          : std_logic_vector(0 to LANE_DATA_WIDTH-1)     := X"0000000000000000";
  signal r_rx_src_ready     : std_logic                                    := '0';
  signal data_err_count_r   : std_logic_vector (0 to 8-1);
  signal pdu_lfsr_r         : std_logic_vector(0 to 15)                    := X"0000";
  signal pdu_cmp_data_w     : std_logic_vector(LANE_DATA_WIDTH-1 downto 0) := X"0000000000000000";
  signal pdu_cmp_data_w_r   : std_logic_vector(0 to LANE_DATA_WIDTH-1)     := X"0000000000000000";

begin

--reset_i <= RESET or not(CHANNEL_UP);
  reset_i <= RESET;



  gen_tdata : for a in 0 to STRB_WIDTH-1 generate

    AXIS_UI_RX_TDATA_i(((STRB_WIDTH-1-a)*8) to ((STRB_WIDTH-1-a)*8)+7) <= AXIS_UI_RX_TDATA(((STRB_WIDTH-1-a)*8)+7 downto ((STRB_WIDTH-1-a)*8));
  end generate gen_tdata;

  process(USER_CLK)
  begin
    if rising_edge(USER_CLK) then
      r_rx_data      <= AXIS_UI_RX_TDATA_i;
      r_rx_src_ready <= not AXIS_UI_RX_TVALID;
    end if;
  end process;
  -----------------------------------------------------------------------------
  --Pseudo data algorithm to generate the same random data as Fram_G
  ----------------------------------------------------------------------------                                      
  process(USER_CLK, reset_i)
  begin
    if reset_i = '1' then
      pdu_lfsr_r <= X"ABCD";            --initial seed to start
    elsif rising_edge(USER_CLK) then
      if (r_rx_src_ready = '0') then
        pdu_lfsr_r <= (not((pdu_lfsr_r(3))xor(pdu_lfsr_r(12))xor(pdu_lfsr_r(14))xor(pdu_lfsr_r(15)))&(pdu_lfsr_r(0 to 14)));
      end if;
    end if;
  end process;

  pdu_cmp_data_w <= pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15)&pdu_lfsr_r(0 to 15);

-------------------------------------------------------------------------------
-- Final data to compare
-------------------------------------------------------------------------------

  pdu_cmp_data_w_r <= pdu_cmp_data_w(63)&pdu_cmp_data_w(62)&pdu_cmp_data_w(61)&pdu_cmp_data_w(60)&
                      pdu_cmp_data_w(59)&pdu_cmp_data_w(58)&pdu_cmp_data_w(57)&pdu_cmp_data_w(56)&
                      pdu_cmp_data_w(55)&pdu_cmp_data_w(54)&pdu_cmp_data_w(53)&pdu_cmp_data_w(52)&
                      pdu_cmp_data_w(51)&pdu_cmp_data_w(50)&pdu_cmp_data_w(49)&pdu_cmp_data_w(48)&
                      pdu_cmp_data_w(47)&pdu_cmp_data_w(46)&pdu_cmp_data_w(45)&pdu_cmp_data_w(44)&
                      pdu_cmp_data_w(43)&pdu_cmp_data_w(42)&pdu_cmp_data_w(41)&pdu_cmp_data_w(40)&
                      pdu_cmp_data_w(39)&pdu_cmp_data_w(38)&pdu_cmp_data_w(37)&pdu_cmp_data_w(36)&
                      pdu_cmp_data_w(35)&pdu_cmp_data_w(34)&pdu_cmp_data_w(33)&pdu_cmp_data_w(32)&
                      pdu_cmp_data_w(31)&pdu_cmp_data_w(30)&pdu_cmp_data_w(29)&pdu_cmp_data_w(28)&
                      pdu_cmp_data_w(27)&pdu_cmp_data_w(26)&pdu_cmp_data_w(25)&pdu_cmp_data_w(24)&
                      pdu_cmp_data_w(23)&pdu_cmp_data_w(22)&pdu_cmp_data_w(21)&pdu_cmp_data_w(20)&
                      pdu_cmp_data_w(19)&pdu_cmp_data_w(18)&pdu_cmp_data_w(17)&pdu_cmp_data_w(16)&
                      pdu_cmp_data_w(15)&pdu_cmp_data_w(14)&pdu_cmp_data_w(13)&pdu_cmp_data_w(12)&
                      pdu_cmp_data_w(11)&pdu_cmp_data_w(10)&pdu_cmp_data_w(9)&pdu_cmp_data_w(8)&
                      pdu_cmp_data_w(7)&pdu_cmp_data_w(6)&pdu_cmp_data_w(5)&pdu_cmp_data_w(4)&
                      pdu_cmp_data_w(3)&pdu_cmp_data_w(2)&pdu_cmp_data_w(1)&pdu_cmp_data_w(0);

-- Data error counter

process(USER_CLK)
begin
	if reset_i ='1' then
		data_err_count_r <=(others=> '0'); 
	elsif rising_edge(USER_CLK) then
	   if r_rx_src_ready='0' then
	    if  data_err_count_r= 255 then
	       data_err_count_r <=(others=> '0'); 
		elsif (pdu_cmp_data_w_r/=r_rx_data ) then
			data_err_count_r <= data_err_count_r + 1;
		end if;
	end if; 
end if;
end process;

DATA_ERR_COUNT<=data_err_count_r;

end architecture rtl;
